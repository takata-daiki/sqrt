library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity bC is
  port( S_BUS_C : inout std_logic_vector(15 downto 0));
end bC;

architecture BEHAVIOR of bC is
begin
end BEHAVIOR;
